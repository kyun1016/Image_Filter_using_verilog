// ../../list_tx_model.f 

package pkg_tx_data;
  `include "cls_read_ppm.sv"
  `include "cls_apb.sv"
endpackage

